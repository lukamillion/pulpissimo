//-----------------------------------------------------------------------------
// Title   : PULPissimo Top
// -----------------------------------------------------------------------------
// File    : pulpissimo.sv
// Author  : Manuel Eggimann <meggimann@iis.ee.ethz.ch>
// Created : 19.04.2022
// -----------------------------------------------------------------------------
// Description :
//
// This is the default toplevel of pulpissimo used as the basis for ASIC
// implementations and RTL simulation. It instantiates the following clock
// generation and pad multiplexing IP as well as the `soc_domain` (which wraps
// almost the entire logic of pulpissimo from the external pulp_soc repository).
// The `pulp_soc` repository is shared between the single core variant
// PULPissimo and the multi-core variant pulp-open.
//
//-----------------------------------------------------------------------------
// Copyright (C) 2022 ETH Zurich, University of Bologna Copyright and related
// rights are licensed under the Solderpad Hardware License, Version 0.51 (the
// "License"); you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law or
// agreed to in writing, software, hardware and materials distributed under this
// License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS
// OF ANY KIND, either express or implied. See the License for the specific
// language governing permissions and limitations under the License.
// SPDX-License-Identifier: SHL-0.51
// -----------------------------------------------------------------------------

module pulpissimo #(
    parameter CORE_TYPE     = 0, // TODO check if still up-to date 0 for RISCY, 1 for IBEX RV32IMC (formerly ZERORISCY), 2 for IBEX RV32EC (formerly MICRORISCY)
    parameter USE_FPU       = 1,
    parameter USE_ZFINX     = 1,
    parameter USE_HWPE      = 0,
    parameter SIM_STDOUT    = 0,
    localparam IO_PAD_COUNT = 32 // Check the README on how to modify the pad count
)(
  // Some platforms (e.g. Verilator) require to feed the clock externally. With
  // the EXTERNAL_CLOCK define we remove all internall clock generation logic.
`ifdef EXTERNAL_CLOCK
  input logic ext_slow_clk_i,
  input logic ext_soc_clk_i,
  input logic ext_per_clk_i,
`else
   // Reference clock for clock internal clock generation
  inout wire pad_refclk_in,
`endif
  // Active-low Asynchronous hard-reset
  inout wire pad_reset_n,
  // Clock Bypass enable. If asserted (active-high) peripheral and soc clock
  // domain will be driven directly by pad_refclk_in (or verilator_slow_clk_i if
  // in built for VERILATOR).
  inout wire pad_clk_byp_en,
  // Boot mode selection. Check bootcode repository for mapping of bootsel
  // values to actual boot mode.
  inout wire pad_bootsel0,
  inout wire pad_bootsel1,
  // JTAG in-system debug interface
  inout wire pad_jtag_tck,
  inout wire pad_jtag_tdi,
  inout wire pad_jtag_tdo,
  inout wire pad_jtag_tms,
  inout wire pad_jtag_trst
  // general purpose pads (since PULPissimo v8.0 any peripheral (including
  // GPIO) can be mapped to any pad any-to-any muxing. Check the latest
  // README.md on description and how to modify the pad count)
  inout wire [IO_PAD_COUNT-1:0] pad_io
);


  //////////////////////////////
  // Clock & Reset Generation //
  //////////////////////////////
`ifndef EXTERNAL_CLOCK
  clock_gen i_clock_rst_gen(

  );
`else

`endif



  ///////////////////////////////
  // APB Chip Control Demuxing //
  ///////////////////////////////


  /////////////////////////////////////////////////
  // Pad Multiplexer (Auto-generated by Padrick) //
  /////////////////////////////////////////////////


  /////////////////
  // SoC Wrapper //
  /////////////////
  soc_domain #(
    .CORE_TYPE  ( CORE_TYPE  ),
    .USE_FPU    ( USE_FPU    ),
    .USE_ZFINX  ( USE_ZFINX  ),
    .USE_HWPE   ( USE_HWPE   ),
    .SIM_STDOUT ( SIM_STDOUT )
  ) i_soc_domain (
    // TODO
  );



endmodule
